module test_lut_n();
//This is a test-bench for the look-up table.  The point is to make sure that different instances of lut_n can
//reference different lookup tables stored in the (`include-d) file, cornerNclk.v.
//
//Ted Golfinopoulos, 13 Mar 2012


endmodule 

